module bPredictor(input clk,
	input [15:0]pc
	);
	
endmodule